library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity data is port(
	fetch   :  in  std_logic;
	data_out  :  out std_logic_vector(37 downto 0));
end data;

architecture b of data is
	
	signal storage_index : unsigned(5 downto 0) := (others => '0');
	type data_storage is array(0 to 50) of std_logic_vector(37 downto 0);
	constant data : data_storage := (
	"10011010110111011011001001010010001111", 
	"01100111101110011100011000001001111011", 
	"00100111101110010100010000001001110001", 
	"01111110011101010000011000001010010110", 
	"11010101111001010000111000001010010101", 
	"11010101111000010000001101100100110010", 
	"11000110101000011000110000101111000010", 
	"11010101110001101010110000110100100001", 
	"11001010101010010100010000001001111000", 
	"01100011101110010100010000001001110001", 
	"01100111101110010011101110011101101101", 
	"11010111111000010011010001100000011000", 
	"01100111101110010100010000001001110001", 
	"01100111110100100011100100100100011110", 
	"11010101110001101000110000110100100001", 
	"11010101111000010001101101001011000000", 
	"10010000011101000000110000001010010101", 
	"11010101111000010000111000001010010101", 
	"00110001111101001100011000001011110001", 
	"01100111101110010000011001100101010000", 
	"11010101111000010000111000101111001001", 
	"11010101110001101000110000110100100011", 
	"11001011101010100100011000001001111000", 
	"01100111101110010011011111111101101000", 
	"11010101111000010010111000001010010101", 
	"10010111010011010100011000001011110000", 
	"01100111101110010100010000001001110001", 
	"01110011110110001000111000101111000001", 
	"11010101110001101000110000110100101001", 
	"11010101111000010011111100111000101101", 
	"01100111101110010100010000001001110001", 
	"01100111101110010100010000001001110001", 
	"10011011010100101000010100001000010110", 
	"01100011101110010011000000000011101110", 
	"11010101111000010000111000101111001001", 
	"11010101110001101001101110111111010000", 
	"01100111101110111100011000001001111011", 
	"00111011000100110000110000001000010101", 
	"11010101111000010000111010001010010101", 
	"01111001001111011100010000001011110011", 
	"01100111101110010100010000001001010001", 
	"01100111110100100000001001101111101000", 
	"11010101110001101000110000110100100001", 
	"11010101111000010000010100000011100001", 
	"01101111101110010100010000001001110001", 
	"01100111101110010011110010100010010111", 
	"10010111011000110100010000001001111001", 
	"01100111101110010100011000100111101101", 
	"11010101111000010000111000101111001001", 
	"11010101110011101011000100000111001111", 
	"10011110100011010000110000010000001110"
	);
	
begin
	
	process (fetch)
	begin
		if rising_edge(fetch) then
			storage_index <= storage_index + 1;
		end if;
	end process;
	
	data_out <= data(to_integer(storage_index));
end b;
